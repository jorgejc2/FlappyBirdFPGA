/*
 * ECE385-HelperTools/PNG-To-Txt
 * Author: Rishi Thakkar
 *
 */

module  frameRAM
(
		// input [2:0] data_In,
		// // input [18:0] write_address, read_address,
		// input [8:0] write_address, read_address,
		// input we, Clk,
		input [11:0] read_address,
		output logic [2:0] data_Out
		// input [15:0] read_address,
		// output logic [23:0] data_Out
);

// mem has width of 3 bits and a total of 400 addresses
// logic [23:0] mem [0:32767];
logic [2:0] mem [0:2499];
// parameter ADDR_WIDTH = 12;
// parameter DATA_WIDTH = 3;
// logic [ADDR_WIDTH-1:0] addr_reg;
initial 
begin
	$readmemh("sprite_bytes/bird.txt",mem);
	// $readmemh("sounds_converted/formatted_sound.txt",mem);
end


// parameter bit [DATA_WIDTH-1:0] mem [0:2**ADDR_WIDTH-1] = '{
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h6,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h4,
// 3'h4,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h4,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h5,
// 3'h2,
// 3'h1,
// 3'h1,
// 3'h1,
// 3'h4,
// 3'h4,
// 3'h2,
// 3'h5,
// 3'h3,
// 3'h4,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h5,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h3,
// 3'h5,
// 3'h2
// };

// initial
// begin
// 	 $readmemh("sprite_bytes/bird.txt", mem);
// end


// always_ff @ (posedge Clk) begin
// 	if (we)
// 		mem[write_address] <= data_In;
// 	data_Out<= mem[read_address];
// end

assign data_Out = mem[read_address];

endmodule
