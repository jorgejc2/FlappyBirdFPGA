//-------------------------------------------------------------------------
//                                                                       --
//                                                                       --
//      For use with ECE 385 Lab 62                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab62 (

      ///////// Clocks /////////
      input     MAX10_CLK1_50, 

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,


      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);




logic Reset_h, vssig, blank, sync, VGA_Clk;


//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
	logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
	logic [1:0] signs;
	logic [1:0] hundreds;
	logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig, greenpipe1_x, greenpipe1_y,greenpipe2_x, greenpipe2_y,
	greenpipe3_x, greenpipe3_y, greenpipe4_x, greenpipe4_y,
	CLOUD1_x, CLOUD1_y , CLOUD2_x, CLOUD2_y  ,CLOUD3_x ,CLOUD3_y  , CLOUD4_x ,
    CLOUD4_y ,
    CLOUD5_x ,CLOUD5_y;
	logic [7:0] Red, Blue, Green;
	logic [7:0] keycode;
	logic [26:0] score_num;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ; 
	assign USB_IRQ = ARDUINO_IO[9];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[7] = USB_RST;//USB reset 
	assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
	assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt
	
	//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
	assign ARDUINO_IO[6] = 1'b1;
	
	//HEX drivers to convert numbers to HEX output
	HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
	assign HEX4[7] = 1'b1;
	
	HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
	assign HEX3[7] = 1'b1;
	
	HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
	assign HEX1[7] = 1'b1;
	
	HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
	assign HEX0[7] = 1'b1;
	
	//fill in the hundreds digit as well as the negative sign
	assign HEX5 = {1'b1, ~signs[1], 3'b111, ~hundreds[1], ~hundreds[1], 1'b1};
	assign HEX2 = {1'b1, ~signs[0], 3'b111, ~hundreds[0], ~hundreds[0], 1'b1};
	
	
	//Assign one button to reset
	assign {Reset_h}=~ (KEY[0]);

	//Our A/D converter is only 12 bit
	assign VGA_R = Red[7:4];
	assign VGA_B = Blue[7:4];
	assign VGA_G = Green[7:4];
	
	
	lab62soc u0 (
		.clk_clk                           (MAX10_CLK1_50),  //clk.clk
		.reset_reset_n                     (1'b1),           //reset.reset_n
		.altpll_0_locked_conduit_export    (),               //altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (),               //altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),               //altpll_0_areset_conduit.export
		.key_external_connection_export    (KEY),            //key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),                            //clk_sdram.clk
		.sdram_wire_addr(DRAM_ADDR),                         //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                             //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),                       //.cas_n
		.sdram_wire_cke(DRAM_CKE),                           //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                         //.cs_n
		.sdram_wire_dq(DRAM_DQ),                             //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),              //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),                       //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                         //.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.hex_digits_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),
		// .leds_export({hundreds, signs, LEDR}),
		.keycode_export(keycode)
		
	 );

logic [9:0] x1, y1, x2, y2, x3, x4, x5;
    assign x1 = 50;
    assign y1 = 200;
	assign y2 = 100;
    assign x2 = 200;
    assign x3 = 350;
    assign x4 = 500;
    assign x5 = 600;
//instantiate a vga_controller, ball, and color_mapper here with the ports.

ball ball0 (.Reset(Reset_h), .frame_clk(VGA_VS),.keycode(keycode),.BallX(ballxsig), .BallY(ballysig), .BallS(ballsizesig) );

vga_controller vga0( .Clk(MAX10_CLK1_50), .Reset(Reset_h),.hs(VGA_HS), 
								              .vs(VGA_VS),
												  .pixel_clk(VGA_Clk), 
												  .blank(blank),     
												  .sync(sync), .DrawX(drawxsig),     
								              .DrawY(drawysig) );

color_mapper color0(.Clk(MAX10_CLK1_50), .Reset(Reset_h), .VGA_Clk(VGA_VS), .Blank(blank), .BallX(ballxsig), .BallY(ballysig), .DrawX(drawxsig), .DrawY(drawysig), .Ball_size(ballsizesig),
							.Red(Red), .Green(Green), .Blue(Blue), .eightOut(LEDR[7:0]), .keycode(keycode), 
							.pipe1X(greenpipe1_x), .pipe1Y(greenpipe1_y), .pipe2X(greenpipe2_x), .pipe2Y(greenpipe2_y),
							.pipe3X(greenpipe3_x), .pipe3Y(greenpipe3_y), .pipe4X(greenpipe4_x), .pipe4Y(greenpipe4_y), 
							.cloud1X(CLOUD1_x), .cloud1Y(CLOUD1_y), 
							.cloud2X(CLOUD2_x), .cloud2Y(CLOUD2_y), 
							.cloud3X(CLOUD3_x), .cloud3Y(CLOUD3_y), 
							.cloud4X(CLOUD4_x), .cloud4Y(CLOUD4_y), 
							.cloud5X(CLOUD5_x), .cloud5Y(CLOUD5_y),  .score(score_num)
							);

greenpipe1 greenpipe1_0 (.Reset(Reset_h), .frame_clk(VGA_VS),.keycode(8'h04),.BallX(greenpipe1_x),
    .BallY(greenpipe1_y), .BallS(), .score(score_num));
greenpipe2 greenpipe2_0 (.Reset(Reset_h), .frame_clk(VGA_VS),.keycode(8'h04),.BallX(greenpipe2_x),
.BallY(greenpipe2_y), .BallS() , .score(score_num));
greenpipe3 greenpipe3_0 (.Reset(Reset_h), .frame_clk(VGA_VS),.keycode(8'h04),.BallX(greenpipe3_x),
.BallY(greenpipe3_y), .BallS() , .score(score_num));
greenpipe4 greenpipe4_0 (.Reset(Reset_h), .frame_clk(VGA_VS),.keycode(8'h04),.BallX(greenpipe4_x),
    .BallY(greenpipe4_y), .BallS(), .score(score_num));

cloudMovements cloudMovements1(.Reset(Reset_h), .frame_clk(VGA_VS),
               .BallX(CLOUD1_x), .BallY(CLOUD1_y), .BallS(), .startX(x1), .startY(y1), .keycode(8'h04) );
    cloudMovements cloudMovements2(.Reset(Reset_h), .frame_clk(VGA_VS),
               .BallX(CLOUD2_x), .BallY(CLOUD2_y), .BallS(), .startX(x2), .startY(y2), .keycode(8'h04) );
    cloudMovements cloudMovements3(.Reset(Reset_h), .frame_clk(VGA_VS),
               .BallX(CLOUD3_x), .BallY(CLOUD3_y), .BallS(), .startX(x3), .startY(y1), .keycode(8'h04) );
    cloudMovements cloudMovements4(.Reset(Reset_h), .frame_clk(VGA_VS),
               .BallX(CLOUD4_x), .BallY(CLOUD4_y), .BallS(), .startX(x4), .startY(y2), .keycode(8'h04) );
    cloudMovements cloudMovements5(.Reset(Reset_h), .frame_clk(VGA_VS),
               .BallX(CLOUD5_x), .BallY(CLOUD5_y), .BallS(), .startX(x5), .startY(y1), .keycode(8'h04) );

endmodule
